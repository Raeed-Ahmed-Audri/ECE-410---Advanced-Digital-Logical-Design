----------------------------------------------------------------------------------
-- Filename : mux_tb.vhdl
-- Author : Antonio Alejandro Andara Lara
-- Date : 31-Oct-2023
-- Design Name: mux_tb
-- Project Name: ECE 410 lab 3 2023
-- Description : testbench for the multiplexer of the simple CPU design
-- Revision 1.01 - File Modified by Antonio Andara (October 28, 2024)
-- Additional Comments:
-- Copyright : University of Alberta, 2023
-- License : CC0 1.0 Universal
----------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mux4_tb IS
END mux4_tb;

ARCHITECTURE sim OF mux4_tb IS

    SIGNAL in0    : STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in1    : STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in2    : STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL in3    : STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL mux_sel : STD_LOGIC_VECTOR(1 DOWNTO 0)  := "00";
    SIGNAL mux_out : STD_LOGIC_VECTOR(15 DOWNTO 0);

BEGIN
    -- Instantiate the Unit Under Test (UUT)

    uut : ENTITY work.mux4(Dataflow)
        PORT MAP(
            in0 => in0,
            in1 => in1,
            in2 => in2,
            in3 => in3,
            mux_sel => mux_sel,
            mux_out => mux_out           
        );

    stimulus : PROCESS
    BEGIN
        -- Setup test data
        in0     <= "1010101010101010"; --16 bits wide
        in1     <= "1100110011001100";
        in2     <= "1111000011110000";
        in3     <= "0000111100001111";

        -- Select in0
        mux_sel <= "00";
        WAIT FOR 20 ns;

        -- Assertion to check if output matches in0
        ASSERT (mux_out = in0)
        REPORT "Mismatch for mux_sel = 00!"
            SEVERITY ERROR;
            
           -- Select in1
        mux_sel <= "01";
        WAIT FOR 20 ns;

        -- Assertion to check if output matches in1
        ASSERT (mux_out = in1)
        REPORT "Mismatch for mux_sel = 01!"
            SEVERITY ERROR;
            
           -- Select in2
        mux_sel <= "10";
        WAIT FOR 20 ns;

        -- Assertion to check if output matches in2
        ASSERT (mux_out = in2)
        REPORT "Mismatch for mux_sel = 10!"
            SEVERITY ERROR;
            
          -- Select in3
        mux_sel <= "11";
        WAIT FOR 20 ns;

        -- Assertion to check if output matches in3
        ASSERT (mux_out = in3)
        REPORT "Mismatch for mux_sel = 11!"
            SEVERITY ERROR;

        -- End the test
        WAIT;
    END PROCESS stimulus;

END sim;
